`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.06.2025 18:45:28
// Design Name: 
// Module Name: cos_lut
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cos_lut (
    input wire [15:0] phase,             // 16-bit phase accumulator
    output reg signed [15:0] cos_val     // 16-bit signed cosine output
);

    // Use the top 10 bits to index into 1024-entry LUT
    wire [9:0] addr = phase[15:6];

    // Cosine lookup table (scaled by 16384 for Q1.14 format)
    reg signed [15:0] lut [0:1023];

    initial begin
    lut[0] = 16'sd16384;
    lut[1] = 16'sd16384;
    lut[2] = 16'sd16383;
    lut[3] = 16'sd16381;
    lut[4] = 16'sd16379;
    lut[5] = 16'sd16376;
    lut[6] = 16'sd16373;
    lut[7] = 16'sd16369;
    lut[8] = 16'sd16364;
    lut[9] = 16'sd16359;
    lut[10] = 16'sd16353;
    lut[11] = 16'sd16347;
    lut[12] = 16'sd16340;
    lut[13] = 16'sd16332;
    lut[14] = 16'sd16324;
    lut[15] = 16'sd16315;
    lut[16] = 16'sd16305;
    lut[17] = 16'sd16295;
    lut[18] = 16'sd16284;
    lut[19] = 16'sd16273;
    lut[20] = 16'sd16261;
    lut[21] = 16'sd16248;
    lut[22] = 16'sd16235;
    lut[23] = 16'sd16221;
    lut[24] = 16'sd16207;
    lut[25] = 16'sd16192;
    lut[26] = 16'sd16176;
    lut[27] = 16'sd16160;
    lut[28] = 16'sd16143;
    lut[29] = 16'sd16125;
    lut[30] = 16'sd16107;
    lut[31] = 16'sd16088;
    lut[32] = 16'sd16069;
    lut[33] = 16'sd16049;
    lut[34] = 16'sd16029;
    lut[35] = 16'sd16008;
    lut[36] = 16'sd15986;
    lut[37] = 16'sd15964;
    lut[38] = 16'sd15941;
    lut[39] = 16'sd15917;
    lut[40] = 16'sd15893;
    lut[41] = 16'sd15868;
    lut[42] = 16'sd15843;
    lut[43] = 16'sd15817;
    lut[44] = 16'sd15791;
    lut[45] = 16'sd15763;
    lut[46] = 16'sd15736;
    lut[47] = 16'sd15707;
    lut[48] = 16'sd15679;
    lut[49] = 16'sd15649;
    lut[50] = 16'sd15619;
    lut[51] = 16'sd15588;
    lut[52] = 16'sd15557;
    lut[53] = 16'sd15525;
    lut[54] = 16'sd15493;
    lut[55] = 16'sd15460;
    lut[56] = 16'sd15426;
    lut[57] = 16'sd15392;
    lut[58] = 16'sd15357;
    lut[59] = 16'sd15322;
    lut[60] = 16'sd15286;
    lut[61] = 16'sd15250;
    lut[62] = 16'sd15213;
    lut[63] = 16'sd15175;
    lut[64] = 16'sd15137;
    lut[65] = 16'sd15098;
    lut[66] = 16'sd15059;
    lut[67] = 16'sd15019;
    lut[68] = 16'sd14978;
    lut[69] = 16'sd14937;
    lut[70] = 16'sd14896;
    lut[71] = 16'sd14854;
    lut[72] = 16'sd14811;
    lut[73] = 16'sd14768;
    lut[74] = 16'sd14724;
    lut[75] = 16'sd14680;
    lut[76] = 16'sd14635;
    lut[77] = 16'sd14589;
    lut[78] = 16'sd14543;
    lut[79] = 16'sd14497;
    lut[80] = 16'sd14449;
    lut[81] = 16'sd14402;
    lut[82] = 16'sd14354;
    lut[83] = 16'sd14305;
    lut[84] = 16'sd14256;
    lut[85] = 16'sd14206;
    lut[86] = 16'sd14155;
    lut[87] = 16'sd14104;
    lut[88] = 16'sd14053;
    lut[89] = 16'sd14001;
    lut[90] = 16'sd13949;
    lut[91] = 16'sd13896;
    lut[92] = 16'sd13842;
    lut[93] = 16'sd13788;
    lut[94] = 16'sd13733;
    lut[95] = 16'sd13678;
    lut[96] = 16'sd13623;
    lut[97] = 16'sd13567;
    lut[98] = 16'sd13510;
    lut[99] = 16'sd13453;
    lut[100] = 16'sd13395;
    lut[101] = 16'sd13337;
    lut[102] = 16'sd13279;
    lut[103] = 16'sd13219;
    lut[104] = 16'sd13160;
    lut[105] = 16'sd13100;
    lut[106] = 16'sd13039;
    lut[107] = 16'sd12978;
    lut[108] = 16'sd12916;
    lut[109] = 16'sd12854;
    lut[110] = 16'sd12792;
    lut[111] = 16'sd12729;
    lut[112] = 16'sd12665;
    lut[113] = 16'sd12601;
    lut[114] = 16'sd12537;
    lut[115] = 16'sd12472;
    lut[116] = 16'sd12406;
    lut[117] = 16'sd12340;
    lut[118] = 16'sd12274;
    lut[119] = 16'sd12207;
    lut[120] = 16'sd12140;
    lut[121] = 16'sd12072;
    lut[122] = 16'sd12004;
    lut[123] = 16'sd11935;
    lut[124] = 16'sd11866;
    lut[125] = 16'sd11797;
    lut[126] = 16'sd11727;
    lut[127] = 16'sd11656;
    lut[128] = 16'sd11585;
    lut[129] = 16'sd11514;
    lut[130] = 16'sd11442;
    lut[131] = 16'sd11370;
    lut[132] = 16'sd11297;
    lut[133] = 16'sd11224;
    lut[134] = 16'sd11151;
    lut[135] = 16'sd11077;
    lut[136] = 16'sd11003;
    lut[137] = 16'sd10928;
    lut[138] = 16'sd10853;
    lut[139] = 16'sd10778;
    lut[140] = 16'sd10702;
    lut[141] = 16'sd10625;
    lut[142] = 16'sd10549;
    lut[143] = 16'sd10471;
    lut[144] = 16'sd10394;
    lut[145] = 16'sd10316;
    lut[146] = 16'sd10238;
    lut[147] = 16'sd10159;
    lut[148] = 16'sd10080;
    lut[149] = 16'sd10001;
    lut[150] = 16'sd9921;
    lut[151] = 16'sd9841;
    lut[152] = 16'sd9760;
    lut[153] = 16'sd9679;
    lut[154] = 16'sd9598;
    lut[155] = 16'sd9516;
    lut[156] = 16'sd9434;
    lut[157] = 16'sd9352;
    lut[158] = 16'sd9269;
    lut[159] = 16'sd9186;
    lut[160] = 16'sd9102;
    lut[161] = 16'sd9019;
    lut[162] = 16'sd8935;
    lut[163] = 16'sd8850;
    lut[164] = 16'sd8765;
    lut[165] = 16'sd8680;
    lut[166] = 16'sd8595;
    lut[167] = 16'sd8509;
    lut[168] = 16'sd8423;
    lut[169] = 16'sd8337;
    lut[170] = 16'sd8250;
    lut[171] = 16'sd8163;
    lut[172] = 16'sd8076;
    lut[173] = 16'sd7988;
    lut[174] = 16'sd7900;
    lut[175] = 16'sd7812;
    lut[176] = 16'sd7723;
    lut[177] = 16'sd7635;
    lut[178] = 16'sd7545;
    lut[179] = 16'sd7456;
    lut[180] = 16'sd7366;
    lut[181] = 16'sd7276;
    lut[182] = 16'sd7186;
    lut[183] = 16'sd7096;
    lut[184] = 16'sd7005;
    lut[185] = 16'sd6914;
    lut[186] = 16'sd6823;
    lut[187] = 16'sd6731;
    lut[188] = 16'sd6639;
    lut[189] = 16'sd6547;
    lut[190] = 16'sd6455;
    lut[191] = 16'sd6363;
    lut[192] = 16'sd6270;
    lut[193] = 16'sd6177;
    lut[194] = 16'sd6084;
    lut[195] = 16'sd5990;
    lut[196] = 16'sd5897;
    lut[197] = 16'sd5803;
    lut[198] = 16'sd5708;
    lut[199] = 16'sd5614;
    lut[200] = 16'sd5520;
    lut[201] = 16'sd5425;
    lut[202] = 16'sd5330;
    lut[203] = 16'sd5235;
    lut[204] = 16'sd5139;
    lut[205] = 16'sd5044;
    lut[206] = 16'sd4948;
    lut[207] = 16'sd4852;
    lut[208] = 16'sd4756;
    lut[209] = 16'sd4660;
    lut[210] = 16'sd4563;
    lut[211] = 16'sd4467;
    lut[212] = 16'sd4370;
    lut[213] = 16'sd4273;
    lut[214] = 16'sd4176;
    lut[215] = 16'sd4078;
    lut[216] = 16'sd3981;
    lut[217] = 16'sd3883;
    lut[218] = 16'sd3786;
    lut[219] = 16'sd3688;
    lut[220] = 16'sd3590;
    lut[221] = 16'sd3492;
    lut[222] = 16'sd3393;
    lut[223] = 16'sd3295;
    lut[224] = 16'sd3196;
    lut[225] = 16'sd3098;
    lut[226] = 16'sd2999;
    lut[227] = 16'sd2900;
    lut[228] = 16'sd2801;
    lut[229] = 16'sd2702;
    lut[230] = 16'sd2603;
    lut[231] = 16'sd2503;
    lut[232] = 16'sd2404;
    lut[233] = 16'sd2305;
    lut[234] = 16'sd2205;
    lut[235] = 16'sd2105;
    lut[236] = 16'sd2006;
    lut[237] = 16'sd1906;
    lut[238] = 16'sd1806;
    lut[239] = 16'sd1706;
    lut[240] = 16'sd1606;
    lut[241] = 16'sd1506;
    lut[242] = 16'sd1406;
    lut[243] = 16'sd1306;
    lut[244] = 16'sd1205;
    lut[245] = 16'sd1105;
    lut[246] = 16'sd1005;
    lut[247] = 16'sd904;
    lut[248] = 16'sd804;
    lut[249] = 16'sd704;
    lut[250] = 16'sd603;
    lut[251] = 16'sd503;
    lut[252] = 16'sd402;
    lut[253] = 16'sd302;
    lut[254] = 16'sd201;
    lut[255] = 16'sd101;
    lut[256] = 16'sd0;
    lut[257] = -16'sd101;
    lut[258] = -16'sd201;
    lut[259] = -16'sd302;
    lut[260] = -16'sd402;
    lut[261] = -16'sd503;
    lut[262] = -16'sd603;
    lut[263] = -16'sd704;
    lut[264] = -16'sd804;
    lut[265] = -16'sd904;
    lut[266] = -16'sd1005;
    lut[267] = -16'sd1105;
    lut[268] = -16'sd1205;
    lut[269] = -16'sd1306;
    lut[270] = -16'sd1406;
    lut[271] = -16'sd1506;
    lut[272] = -16'sd1606;
    lut[273] = -16'sd1706;
    lut[274] = -16'sd1806;
    lut[275] = -16'sd1906;
    lut[276] = -16'sd2006;
    lut[277] = -16'sd2105;
    lut[278] = -16'sd2205;
    lut[279] = -16'sd2305;
    lut[280] = -16'sd2404;
    lut[281] = -16'sd2503;
    lut[282] = -16'sd2603;
    lut[283] = -16'sd2702;
    lut[284] = -16'sd2801;
    lut[285] = -16'sd2900;
    lut[286] = -16'sd2999;
    lut[287] = -16'sd3098;
    lut[288] = -16'sd3196;
    lut[289] = -16'sd3295;
    lut[290] = -16'sd3393;
    lut[291] = -16'sd3492;
    lut[292] = -16'sd3590;
    lut[293] = -16'sd3688;
    lut[294] = -16'sd3786;
    lut[295] = -16'sd3883;
    lut[296] = -16'sd3981;
    lut[297] = -16'sd4078;
    lut[298] = -16'sd4176;
    lut[299] = -16'sd4273;
    lut[300] = -16'sd4370;
    lut[301] = -16'sd4467;
    lut[302] = -16'sd4563;
    lut[303] = -16'sd4660;
    lut[304] = -16'sd4756;
    lut[305] = -16'sd4852;
    lut[306] = -16'sd4948;
    lut[307] = -16'sd5044;
    lut[308] = -16'sd5139;
    lut[309] = -16'sd5235;
    lut[310] = -16'sd5330;
    lut[311] = -16'sd5425;
    lut[312] = -16'sd5520;
    lut[313] = -16'sd5614;
    lut[314] = -16'sd5708;
    lut[315] = -16'sd5803;
    lut[316] = -16'sd5897;
    lut[317] = -16'sd5990;
    lut[318] = -16'sd6084;
    lut[319] = -16'sd6177;
    lut[320] = -16'sd6270;
    lut[321] = -16'sd6363;
    lut[322] = -16'sd6455;
    lut[323] = -16'sd6547;
    lut[324] = -16'sd6639;
    lut[325] = -16'sd6731;
    lut[326] = -16'sd6823;
    lut[327] = -16'sd6914;
    lut[328] = -16'sd7005;
    lut[329] = -16'sd7096;
    lut[330] = -16'sd7186;
    lut[331] = -16'sd7276;
    lut[332] = -16'sd7366;
    lut[333] = -16'sd7456;
    lut[334] = -16'sd7545;
    lut[335] = -16'sd7635;
    lut[336] = -16'sd7723;
    lut[337] = -16'sd7812;
    lut[338] = -16'sd7900;
    lut[339] = -16'sd7988;
    lut[340] = -16'sd8076;
    lut[341] = -16'sd8163;
    lut[342] = -16'sd8250;
    lut[343] = -16'sd8337;
    lut[344] = -16'sd8423;
    lut[345] = -16'sd8509;
    lut[346] = -16'sd8595;
    lut[347] = -16'sd8680;
    lut[348] = -16'sd8765;
    lut[349] = -16'sd8850;
    lut[350] = -16'sd8935;
    lut[351] = -16'sd9019;
    lut[352] = -16'sd9102;
    lut[353] = -16'sd9186;
    lut[354] = -16'sd9269;
    lut[355] = -16'sd9352;
    lut[356] = -16'sd9434;
    lut[357] = -16'sd9516;
    lut[358] = -16'sd9598;
    lut[359] = -16'sd9679;
    lut[360] = -16'sd9760;
    lut[361] = -16'sd9841;
    lut[362] = -16'sd9921;
    lut[363] = -16'sd10001;
    lut[364] = -16'sd10080;
    lut[365] = -16'sd10159;
    lut[366] = -16'sd10238;
    lut[367] = -16'sd10316;
    lut[368] = -16'sd10394;
    lut[369] = -16'sd10471;
    lut[370] = -16'sd10549;
    lut[371] = -16'sd10625;
    lut[372] = -16'sd10702;
    lut[373] = -16'sd10778;
    lut[374] = -16'sd10853;
    lut[375] = -16'sd10928;
    lut[376] = -16'sd11003;
    lut[377] = -16'sd11077;
    lut[378] = -16'sd11151;
    lut[379] = -16'sd11224;
    lut[380] = -16'sd11297;
    lut[381] = -16'sd11370;
    lut[382] = -16'sd11442;
    lut[383] = -16'sd11514;
    lut[384] = -16'sd11585;
    lut[385] = -16'sd11656;
    lut[386] = -16'sd11727;
    lut[387] = -16'sd11797;
    lut[388] = -16'sd11866;
    lut[389] = -16'sd11935;
    lut[390] = -16'sd12004;
    lut[391] = -16'sd12072;
    lut[392] = -16'sd12140;
    lut[393] = -16'sd12207;
    lut[394] = -16'sd12274;
    lut[395] = -16'sd12340;
    lut[396] = -16'sd12406;
    lut[397] = -16'sd12472;
    lut[398] = -16'sd12537;
    lut[399] = -16'sd12601;
    lut[400] = -16'sd12665;
    lut[401] = -16'sd12729;
    lut[402] = -16'sd12792;
    lut[403] = -16'sd12854;
    lut[404] = -16'sd12916;
    lut[405] = -16'sd12978;
    lut[406] = -16'sd13039;
    lut[407] = -16'sd13100;
    lut[408] = -16'sd13160;
    lut[409] = -16'sd13219;
    lut[410] = -16'sd13279;
    lut[411] = -16'sd13337;
    lut[412] = -16'sd13395;
    lut[413] = -16'sd13453;
    lut[414] = -16'sd13510;
    lut[415] = -16'sd13567;
    lut[416] = -16'sd13623;
    lut[417] = -16'sd13678;
    lut[418] = -16'sd13733;
    lut[419] = -16'sd13788;
    lut[420] = -16'sd13842;
    lut[421] = -16'sd13896;
    lut[422] = -16'sd13949;
    lut[423] = -16'sd14001;
    lut[424] = -16'sd14053;
    lut[425] = -16'sd14104;
    lut[426] = -16'sd14155;
    lut[427] = -16'sd14206;
    lut[428] = -16'sd14256;
    lut[429] = -16'sd14305;
    lut[430] = -16'sd14354;
    lut[431] = -16'sd14402;
    lut[432] = -16'sd14449;
    lut[433] = -16'sd14497;
    lut[434] = -16'sd14543;
    lut[435] = -16'sd14589;
    lut[436] = -16'sd14635;
    lut[437] = -16'sd14680;
    lut[438] = -16'sd14724;
    lut[439] = -16'sd14768;
    lut[440] = -16'sd14811;
    lut[441] = -16'sd14854;
    lut[442] = -16'sd14896;
    lut[443] = -16'sd14937;
    lut[444] = -16'sd14978;
    lut[445] = -16'sd15019;
    lut[446] = -16'sd15059;
    lut[447] = -16'sd15098;
    lut[448] = -16'sd15137;
    lut[449] = -16'sd15175;
    lut[450] = -16'sd15213;
    lut[451] = -16'sd15250;
    lut[452] = -16'sd15286;
    lut[453] = -16'sd15322;
    lut[454] = -16'sd15357;
    lut[455] = -16'sd15392;
    lut[456] = -16'sd15426;
    lut[457] = -16'sd15460;
    lut[458] = -16'sd15493;
    lut[459] = -16'sd15525;
    lut[460] = -16'sd15557;
    lut[461] = -16'sd15588;
    lut[462] = -16'sd15619;
    lut[463] = -16'sd15649;
    lut[464] = -16'sd15679;
    lut[465] = -16'sd15707;
    lut[466] = -16'sd15736;
    lut[467] = -16'sd15763;
    lut[468] = -16'sd15791;
    lut[469] = -16'sd15817;
    lut[470] = -16'sd15843;
    lut[471] = -16'sd15868;
    lut[472] = -16'sd15893;
    lut[473] = -16'sd15917;
    lut[474] = -16'sd15941;
    lut[475] = -16'sd15964;
    lut[476] = -16'sd15986;
    lut[477] = -16'sd16008;
    lut[478] = -16'sd16029;
    lut[479] = -16'sd16049;
    lut[480] = -16'sd16069;
    lut[481] = -16'sd16088;
    lut[482] = -16'sd16107;
    lut[483] = -16'sd16125;
    lut[484] = -16'sd16143;
    lut[485] = -16'sd16160;
    lut[486] = -16'sd16176;
    lut[487] = -16'sd16192;
    lut[488] = -16'sd16207;
    lut[489] = -16'sd16221;
    lut[490] = -16'sd16235;
    lut[491] = -16'sd16248;
    lut[492] = -16'sd16261;
    lut[493] = -16'sd16273;
    lut[494] = -16'sd16284;
    lut[495] = -16'sd16295;
    lut[496] = -16'sd16305;
    lut[497] = -16'sd16315;
    lut[498] = -16'sd16324;
    lut[499] = -16'sd16332;
    lut[500] = -16'sd16340;
    lut[501] = -16'sd16347;
    lut[502] = -16'sd16353;
    lut[503] = -16'sd16359;
    lut[504] = -16'sd16364;
    lut[505] = -16'sd16369;
    lut[506] = -16'sd16373;
    lut[507] = -16'sd16376;
    lut[508] = -16'sd16379;
    lut[509] = -16'sd16381;
    lut[510] = -16'sd16383;
    lut[511] = -16'sd16384;
    lut[512] = -16'sd16384;
    lut[513] = -16'sd16384;
    lut[514] = -16'sd16383;
    lut[515] = -16'sd16381;
    lut[516] = -16'sd16379;
    lut[517] = -16'sd16376;
    lut[518] = -16'sd16373;
    lut[519] = -16'sd16369;
    lut[520] = -16'sd16364;
    lut[521] = -16'sd16359;
    lut[522] = -16'sd16353;
    lut[523] = -16'sd16347;
    lut[524] = -16'sd16340;
    lut[525] = -16'sd16332;
    lut[526] = -16'sd16324;
    lut[527] = -16'sd16315;
    lut[528] = -16'sd16305;
    lut[529] = -16'sd16295;
    lut[530] = -16'sd16284;
    lut[531] = -16'sd16273;
    lut[532] = -16'sd16261;
    lut[533] = -16'sd16248;
    lut[534] = -16'sd16235;
    lut[535] = -16'sd16221;
    lut[536] = -16'sd16207;
    lut[537] = -16'sd16192;
    lut[538] = -16'sd16176;
    lut[539] = -16'sd16160;
    lut[540] = -16'sd16143;
    lut[541] = -16'sd16125;
    lut[542] = -16'sd16107;
    lut[543] = -16'sd16088;
    lut[544] = -16'sd16069;
    lut[545] = -16'sd16049;
    lut[546] = -16'sd16029;
    lut[547] = -16'sd16008;
    lut[548] = -16'sd15986;
    lut[549] = -16'sd15964;
    lut[550] = -16'sd15941;
    lut[551] = -16'sd15917;
    lut[552] = -16'sd15893;
    lut[553] = -16'sd15868;
    lut[554] = -16'sd15843;
    lut[555] = -16'sd15817;
    lut[556] = -16'sd15791;
    lut[557] = -16'sd15763;
    lut[558] = -16'sd15736;
    lut[559] = -16'sd15707;
    lut[560] = -16'sd15679;
    lut[561] = -16'sd15649;
    lut[562] = -16'sd15619;
    lut[563] = -16'sd15588;
    lut[564] = -16'sd15557;
    lut[565] = -16'sd15525;
    lut[566] = -16'sd15493;
    lut[567] = -16'sd15460;
    lut[568] = -16'sd15426;
    lut[569] = -16'sd15392;
    lut[570] = -16'sd15357;
    lut[571] = -16'sd15322;
    lut[572] = -16'sd15286;
    lut[573] = -16'sd15250;
    lut[574] = -16'sd15213;
    lut[575] = -16'sd15175;
    lut[576] = -16'sd15137;
    lut[577] = -16'sd15098;
    lut[578] = -16'sd15059;
    lut[579] = -16'sd15019;
    lut[580] = -16'sd14978;
    lut[581] = -16'sd14937;
    lut[582] = -16'sd14896;
    lut[583] = -16'sd14854;
    lut[584] = -16'sd14811;
    lut[585] = -16'sd14768;
    lut[586] = -16'sd14724;
    lut[587] = -16'sd14680;
    lut[588] = -16'sd14635;
    lut[589] = -16'sd14589;
    lut[590] = -16'sd14543;
    lut[591] = -16'sd14497;
    lut[592] = -16'sd14449;
    lut[593] = -16'sd14402;
    lut[594] = -16'sd14354;
    lut[595] = -16'sd14305;
    lut[596] = -16'sd14256;
    lut[597] = -16'sd14206;
    lut[598] = -16'sd14155;
    lut[599] = -16'sd14104;
    lut[600] = -16'sd14053;
    lut[601] = -16'sd14001;
    lut[602] = -16'sd13949;
    lut[603] = -16'sd13896;
    lut[604] = -16'sd13842;
    lut[605] = -16'sd13788;
    lut[606] = -16'sd13733;
    lut[607] = -16'sd13678;
    lut[608] = -16'sd13623;
    lut[609] = -16'sd13567;
    lut[610] = -16'sd13510;
    lut[611] = -16'sd13453;
    lut[612] = -16'sd13395;
    lut[613] = -16'sd13337;
    lut[614] = -16'sd13279;
    lut[615] = -16'sd13219;
    lut[616] = -16'sd13160;
    lut[617] = -16'sd13100;
    lut[618] = -16'sd13039;
    lut[619] = -16'sd12978;
    lut[620] = -16'sd12916;
    lut[621] = -16'sd12854;
    lut[622] = -16'sd12792;
    lut[623] = -16'sd12729;
    lut[624] = -16'sd12665;
    lut[625] = -16'sd12601;
    lut[626] = -16'sd12537;
    lut[627] = -16'sd12472;
    lut[628] = -16'sd12406;
    lut[629] = -16'sd12340;
    lut[630] = -16'sd12274;
    lut[631] = -16'sd12207;
    lut[632] = -16'sd12140;
    lut[633] = -16'sd12072;
    lut[634] = -16'sd12004;
    lut[635] = -16'sd11935;
    lut[636] = -16'sd11866;
    lut[637] = -16'sd11797;
    lut[638] = -16'sd11727;
    lut[639] = -16'sd11656;
    lut[640] = -16'sd11585;
    lut[641] = -16'sd11514;
    lut[642] = -16'sd11442;
    lut[643] = -16'sd11370;
    lut[644] = -16'sd11297;
    lut[645] = -16'sd11224;
    lut[646] = -16'sd11151;
    lut[647] = -16'sd11077;
    lut[648] = -16'sd11003;
    lut[649] = -16'sd10928;
    lut[650] = -16'sd10853;
    lut[651] = -16'sd10778;
    lut[652] = -16'sd10702;
    lut[653] = -16'sd10625;
    lut[654] = -16'sd10549;
    lut[655] = -16'sd10471;
    lut[656] = -16'sd10394;
    lut[657] = -16'sd10316;
    lut[658] = -16'sd10238;
    lut[659] = -16'sd10159;
    lut[660] = -16'sd10080;
    lut[661] = -16'sd10001;
    lut[662] = -16'sd9921;
    lut[663] = -16'sd9841;
    lut[664] = -16'sd9760;
    lut[665] = -16'sd9679;
    lut[666] = -16'sd9598;
    lut[667] = -16'sd9516;
    lut[668] = -16'sd9434;
    lut[669] = -16'sd9352;
    lut[670] = -16'sd9269;
    lut[671] = -16'sd9186;
    lut[672] = -16'sd9102;
    lut[673] = -16'sd9019;
    lut[674] = -16'sd8935;
    lut[675] = -16'sd8850;
    lut[676] = -16'sd8765;
    lut[677] = -16'sd8680;
    lut[678] = -16'sd8595;
    lut[679] = -16'sd8509;
    lut[680] = -16'sd8423;
    lut[681] = -16'sd8337;
    lut[682] = -16'sd8250;
    lut[683] = -16'sd8163;
    lut[684] = -16'sd8076;
    lut[685] = -16'sd7988;
    lut[686] = -16'sd7900;
    lut[687] = -16'sd7812;
    lut[688] = -16'sd7723;
    lut[689] = -16'sd7635;
    lut[690] = -16'sd7545;
    lut[691] = -16'sd7456;
    lut[692] = -16'sd7366;
    lut[693] = -16'sd7276;
    lut[694] = -16'sd7186;
    lut[695] = -16'sd7096;
    lut[696] = -16'sd7005;
    lut[697] = -16'sd6914;
    lut[698] = -16'sd6823;
    lut[699] = -16'sd6731;
    lut[700] = -16'sd6639;
    lut[701] = -16'sd6547;
    lut[702] = -16'sd6455;
    lut[703] = -16'sd6363;
    lut[704] = -16'sd6270;
    lut[705] = -16'sd6177;
    lut[706] = -16'sd6084;
    lut[707] = -16'sd5990;
    lut[708] = -16'sd5897;
    lut[709] = -16'sd5803;
    lut[710] = -16'sd5708;
    lut[711] = -16'sd5614;
    lut[712] = -16'sd5520;
    lut[713] = -16'sd5425;
    lut[714] = -16'sd5330;
    lut[715] = -16'sd5235;
    lut[716] = -16'sd5139;
    lut[717] = -16'sd5044;
    lut[718] = -16'sd4948;
    lut[719] = -16'sd4852;
    lut[720] = -16'sd4756;
    lut[721] = -16'sd4660;
    lut[722] = -16'sd4563;
    lut[723] = -16'sd4467;
    lut[724] = -16'sd4370;
    lut[725] = -16'sd4273;
    lut[726] = -16'sd4176;
    lut[727] = -16'sd4078;
    lut[728] = -16'sd3981;
    lut[729] = -16'sd3883;
    lut[730] = -16'sd3786;
    lut[731] = -16'sd3688;
    lut[732] = -16'sd3590;
    lut[733] = -16'sd3492;
    lut[734] = -16'sd3393;
    lut[735] = -16'sd3295;
    lut[736] = -16'sd3196;
    lut[737] = -16'sd3098;
    lut[738] = -16'sd2999;
    lut[739] = -16'sd2900;
    lut[740] = -16'sd2801;
    lut[741] = -16'sd2702;
    lut[742] = -16'sd2603;
    lut[743] = -16'sd2503;
    lut[744] = -16'sd2404;
    lut[745] = -16'sd2305;
    lut[746] = -16'sd2205;
    lut[747] = -16'sd2105;
    lut[748] = -16'sd2006;
    lut[749] = -16'sd1906;
    lut[750] = -16'sd1806;
    lut[751] = -16'sd1706;
    lut[752] = -16'sd1606;
    lut[753] = -16'sd1506;
    lut[754] = -16'sd1406;
    lut[755] = -16'sd1306;
    lut[756] = -16'sd1205;
    lut[757] = -16'sd1105;
    lut[758] = -16'sd1005;
    lut[759] = -16'sd904;
    lut[760] = -16'sd804;
    lut[761] = -16'sd704;
    lut[762] = -16'sd603;
    lut[763] = -16'sd503;
    lut[764] = -16'sd402;
    lut[765] = -16'sd302;
    lut[766] = -16'sd201;
    lut[767] = -16'sd101;
    lut[768] = 16'sd0;
    lut[769] = 16'sd101;
    lut[770] = 16'sd201;
    lut[771] = 16'sd302;
    lut[772] = 16'sd402;
    lut[773] = 16'sd503;
    lut[774] = 16'sd603;
    lut[775] = 16'sd704;
    lut[776] = 16'sd804;
    lut[777] = 16'sd904;
    lut[778] = 16'sd1005;
    lut[779] = 16'sd1105;
    lut[780] = 16'sd1205;
    lut[781] = 16'sd1306;
    lut[782] = 16'sd1406;
    lut[783] = 16'sd1506;
    lut[784] = 16'sd1606;
    lut[785] = 16'sd1706;
    lut[786] = 16'sd1806;
    lut[787] = 16'sd1906;
    lut[788] = 16'sd2006;
    lut[789] = 16'sd2105;
    lut[790] = 16'sd2205;
    lut[791] = 16'sd2305;
    lut[792] = 16'sd2404;
    lut[793] = 16'sd2503;
    lut[794] = 16'sd2603;
    lut[795] = 16'sd2702;
    lut[796] = 16'sd2801;
    lut[797] = 16'sd2900;
    lut[798] = 16'sd2999;
    lut[799] = 16'sd3098;
    lut[800] = 16'sd3196;
    lut[801] = 16'sd3295;
    lut[802] = 16'sd3393;
    lut[803] = 16'sd3492;
    lut[804] = 16'sd3590;
    lut[805] = 16'sd3688;
    lut[806] = 16'sd3786;
    lut[807] = 16'sd3883;
    lut[808] = 16'sd3981;
    lut[809] = 16'sd4078;
    lut[810] = 16'sd4176;
    lut[811] = 16'sd4273;
    lut[812] = 16'sd4370;
    lut[813] = 16'sd4467;
    lut[814] = 16'sd4563;
    lut[815] = 16'sd4660;
    lut[816] = 16'sd4756;
    lut[817] = 16'sd4852;
    lut[818] = 16'sd4948;
    lut[819] = 16'sd5044;
    lut[820] = 16'sd5139;
    lut[821] = 16'sd5235;
    lut[822] = 16'sd5330;
    lut[823] = 16'sd5425;
    lut[824] = 16'sd5520;
    lut[825] = 16'sd5614;
    lut[826] = 16'sd5708;
    lut[827] = 16'sd5803;
    lut[828] = 16'sd5897;
    lut[829] = 16'sd5990;
    lut[830] = 16'sd6084;
    lut[831] = 16'sd6177;
    lut[832] = 16'sd6270;
    lut[833] = 16'sd6363;
    lut[834] = 16'sd6455;
    lut[835] = 16'sd6547;
    lut[836] = 16'sd6639;
    lut[837] = 16'sd6731;
    lut[838] = 16'sd6823;
    lut[839] = 16'sd6914;
    lut[840] = 16'sd7005;
    lut[841] = 16'sd7096;
    lut[842] = 16'sd7186;
    lut[843] = 16'sd7276;
    lut[844] = 16'sd7366;
    lut[845] = 16'sd7456;
    lut[846] = 16'sd7545;
    lut[847] = 16'sd7635;
    lut[848] = 16'sd7723;
    lut[849] = 16'sd7812;
    lut[850] = 16'sd7900;
    lut[851] = 16'sd7988;
    lut[852] = 16'sd8076;
    lut[853] = 16'sd8163;
    lut[854] = 16'sd8250;
    lut[855] = 16'sd8337;
    lut[856] = 16'sd8423;
    lut[857] = 16'sd8509;
    lut[858] = 16'sd8595;
    lut[859] = 16'sd8680;
    lut[860] = 16'sd8765;
    lut[861] = 16'sd8850;
    lut[862] = 16'sd8935;
    lut[863] = 16'sd9019;
    lut[864] = 16'sd9102;
    lut[865] = 16'sd9186;
    lut[866] = 16'sd9269;
    lut[867] = 16'sd9352;
    lut[868] = 16'sd9434;
    lut[869] = 16'sd9516;
    lut[870] = 16'sd9598;
    lut[871] = 16'sd9679;
    lut[872] = 16'sd9760;
    lut[873] = 16'sd9841;
    lut[874] = 16'sd9921;
    lut[875] = 16'sd10001;
    lut[876] = 16'sd10080;
    lut[877] = 16'sd10159;
    lut[878] = 16'sd10238;
    lut[879] = 16'sd10316;
    lut[880] = 16'sd10394;
    lut[881] = 16'sd10471;
    lut[882] = 16'sd10549;
    lut[883] = 16'sd10625;
    lut[884] = 16'sd10702;
    lut[885] = 16'sd10778;
    lut[886] = 16'sd10853;
    lut[887] = 16'sd10928;
    lut[888] = 16'sd11003;
    lut[889] = 16'sd11077;
    lut[890] = 16'sd11151;
    lut[891] = 16'sd11224;
    lut[892] = 16'sd11297;
    lut[893] = 16'sd11370;
    lut[894] = 16'sd11442;
    lut[895] = 16'sd11514;
    lut[896] = 16'sd11585;
    lut[897] = 16'sd11656;
    lut[898] = 16'sd11727;
    lut[899] = 16'sd11797;
    lut[900] = 16'sd11866;
    lut[901] = 16'sd11935;
    lut[902] = 16'sd12004;
    lut[903] = 16'sd12072;
    lut[904] = 16'sd12140;
    lut[905] = 16'sd12207;
    lut[906] = 16'sd12274;
    lut[907] = 16'sd12340;
    lut[908] = 16'sd12406;
    lut[909] = 16'sd12472;
    lut[910] = 16'sd12537;
    lut[911] = 16'sd12601;
    lut[912] = 16'sd12665;
    lut[913] = 16'sd12729;
    lut[914] = 16'sd12792;
    lut[915] = 16'sd12854;
    lut[916] = 16'sd12916;
    lut[917] = 16'sd12978;
    lut[918] = 16'sd13039;
    lut[919] = 16'sd13100;
    lut[920] = 16'sd13160;
    lut[921] = 16'sd13219;
    lut[922] = 16'sd13279;
    lut[923] = 16'sd13337;
    lut[924] = 16'sd13395;
    lut[925] = 16'sd13453;
    lut[926] = 16'sd13510;
    lut[927] = 16'sd13567;
    lut[928] = 16'sd13623;
    lut[929] = 16'sd13678;
    lut[930] = 16'sd13733;
    lut[931] = 16'sd13788;
    lut[932] = 16'sd13842;
    lut[933] = 16'sd13896;
    lut[934] = 16'sd13949;
    lut[935] = 16'sd14001;
    lut[936] = 16'sd14053;
    lut[937] = 16'sd14104;
    lut[938] = 16'sd14155;
    lut[939] = 16'sd14206;
    lut[940] = 16'sd14256;
    lut[941] = 16'sd14305;
    lut[942] = 16'sd14354;
    lut[943] = 16'sd14402;
    lut[944] = 16'sd14449;
    lut[945] = 16'sd14497;
    lut[946] = 16'sd14543;
    lut[947] = 16'sd14589;
    lut[948] = 16'sd14635;
    lut[949] = 16'sd14680;
    lut[950] = 16'sd14724;
    lut[951] = 16'sd14768;
    lut[952] = 16'sd14811;
    lut[953] = 16'sd14854;
    lut[954] = 16'sd14896;
    lut[955] = 16'sd14937;
    lut[956] = 16'sd14978;
    lut[957] = 16'sd15019;
    lut[958] = 16'sd15059;
    lut[959] = 16'sd15098;
    lut[960] = 16'sd15137;
    lut[961] = 16'sd15175;
    lut[962] = 16'sd15213;
    lut[963] = 16'sd15250;
    lut[964] = 16'sd15286;
    lut[965] = 16'sd15322;
    lut[966] = 16'sd15357;
    lut[967] = 16'sd15392;
    lut[968] = 16'sd15426;
    lut[969] = 16'sd15460;
    lut[970] = 16'sd15493;
    lut[971] = 16'sd15525;
    lut[972] = 16'sd15557;
    lut[973] = 16'sd15588;
    lut[974] = 16'sd15619;
    lut[975] = 16'sd15649;
    lut[976] = 16'sd15679;
    lut[977] = 16'sd15707;
    lut[978] = 16'sd15736;
    lut[979] = 16'sd15763;
    lut[980] = 16'sd15791;
    lut[981] = 16'sd15817;
    lut[982] = 16'sd15843;
    lut[983] = 16'sd15868;
    lut[984] = 16'sd15893;
    lut[985] = 16'sd15917;
    lut[986] = 16'sd15941;
    lut[987] = 16'sd15964;
    lut[988] = 16'sd15986;
    lut[989] = 16'sd16008;
    lut[990] = 16'sd16029;
    lut[991] = 16'sd16049;
    lut[992] = 16'sd16069;
    lut[993] = 16'sd16088;
    lut[994] = 16'sd16107;
    lut[995] = 16'sd16125;
    lut[996] = 16'sd16143;
    lut[997] = 16'sd16160;
    lut[998] = 16'sd16176;
    lut[999] = 16'sd16192;
    lut[1000] = 16'sd16207;
    lut[1001] = 16'sd16221;
    lut[1002] = 16'sd16235;
    lut[1003] = 16'sd16248;
    lut[1004] = 16'sd16261;
    lut[1005] = 16'sd16273;
    lut[1006] = 16'sd16284;
    lut[1007] = 16'sd16295;
    lut[1008] = 16'sd16305;
    lut[1009] = 16'sd16315;
    lut[1010] = 16'sd16324;
    lut[1011] = 16'sd16332;
    lut[1012] = 16'sd16340;
    lut[1013] = 16'sd16347;
    lut[1014] = 16'sd16353;
    lut[1015] = 16'sd16359;
    lut[1016] = 16'sd16364;
    lut[1017] = 16'sd16369;
    lut[1018] = 16'sd16373;
    lut[1019] = 16'sd16376;
    lut[1020] = 16'sd16379;
    lut[1021] = 16'sd16381;
    lut[1022] = 16'sd16383;
    lut[1023] = 16'sd16384;
end

    always @(*) begin
        cos_val = lut[addr];
    end

endmodule

